library IEEE;
use IEEE.STD_LOGIC_1164.all;

package utils is
  function MAX (LEFT, RIGHT: INTEGER) return INTEGER;
  function MIN (LEFT, RIGHT: INTEGER) return INTEGER;
END PACKAGE;