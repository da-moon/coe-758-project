package body cache_pkg is

end cache_pkg;
