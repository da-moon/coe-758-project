
library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
package cache_pkg is
TYPE CACHE_MEMORY IS ARRAY (7 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE MAIN_MEMORY IS ARRAY (7 DOWNTO 0, 31 DOWNTO 0) OF std_logic_vector(7 DOWNTO 0);
TYPE STATE IS (READY_STATE, HIT, READ_DATA, WRITE_DATA, IDLE);

FUNCTION GET_TAG(ARG : IN STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR ;
FUNCTION GET_INDEX(ARG : IN STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR ;
FUNCTION GET_OFFSET(ARG : IN STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR ;


end cache_pkg;

package body cache_pkg is
FUNCTION GET_TAG(ARG : IN STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
VARIABLE tag : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
BEGIN
tag := ARG(15 DOWNTO 8);
RETURN tag;
END;
-- -----------------------------------------------------------------------------------------------------------

FUNCTION GET_INDEX(ARG : IN STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
VARIABLE index : STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
BEGIN
index := ARG(7 DOWNTO 5);
RETURN index;
END;
-- -----------------------------------------------------------------------------------------------------------
FUNCTION GET_OFFSET(ARG : IN STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
VARIABLE offset : STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
BEGIN
offset := ARG(4 DOWNTO 0);
RETURN offset;
END;
end cache_pkg;
