
ARCHITECTURE behaviour OF bram IS
  CONSTANT memTypeLength : INTEGER := 2 ** ADDR - 1;
  TYPE MemType IS ARRAY(0 TO memTypeLength) OF STD_LOGIC_VECTOR(DATA - 1 DOWNTO 0);
  IMPURE FUNCTION InitRamFromFile (ARG : IN STRING) RETURN MemType IS
    -- FILE RamFile : text IS IN ARG;
    FILE RamFile : text;
    VARIABLE fstatus : file_open_status;
    VARIABLE RamFileLine : line;
    VARIABLE RAM : MemType;
  BEGIN
    file_open(fstatus, RamFile, ARG, read_mode);
    FOR I IN MemType'RANGE LOOP
      readline (RamFile, RamFileLine);
      hread (RamFileLine, RAM(I)
      );
    END LOOP;
    file_close(RamFile);
    RETURN RAM;
  END InitRamFromFile;
  SIGNAL mem : MemType := InitRamFromFile(RamFileName);
  SIGNAL do : STD_LOGIC_VECTOR(DATA - 1 DOWNTO 0) := (OTHERS => '0');
BEGIN
  PROCESS (clk)
  BEGIN
    IF EDGE = RISING THEN
      CASE MODE IS
        WHEN READ_FIRST => IF rising_edge(clk) THEN
          do <= mem(to_i(adr));
          IF we = '1' THEN
            mem(to_i(adr)) <= din;
          END IF;
      END IF;
      WHEN WRITE_FIRST => IF rising_edge(clk) THEN
      IF we = '1' THEN
        mem(to_i(adr)) <= din;
        do <= din;
      ELSE
        do <= mem(to_i(adr));
      END IF;
    END IF;
    WHEN NO_CHANGE => IF rising_edge(clk) THEN
    IF we = '1' THEN
      mem(to_i(adr)) <= din;
    ELSE
      do <= mem(to_i(adr));
    END IF;
  END IF;
END CASE;
ELSE
CASE MODE IS
  WHEN READ_FIRST => IF falling_edge(clk) THEN
    do <= mem(to_i(adr));
    IF we = '1' THEN
      mem(to_i(adr)) <= din;
    END IF;
END IF;
WHEN WRITE_FIRST => IF falling_edge(clk) THEN
IF we = '1' THEN
  mem(to_i(adr)) <= din;
  do <= din;
ELSE
  do <= mem(to_i(adr));
END IF;
END IF;
WHEN NO_CHANGE => IF falling_edge(clk) THEN
IF we = '1' THEN
  mem(to_i(adr)) <= din;
ELSE
  do <= mem(to_i(adr));
END IF;
END IF;
END CASE;
END IF;
END PROCESS;
--do <= mem(to_i(adr));
dout <= do;
END behaviour;