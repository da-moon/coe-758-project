LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_TEXTIO.ALL;
USE work.cache_pkg.ALL;
USE work.utils_pkg.ALL;
ENTITY bram IS
  GENERIC (
    ADDR : INTEGER := 10;
    DATA : INTEGER := 32;
    EDGE : EdgeType := RISING;
    MODE : MODEType := NO_CHANGE;
    RamFileName : STRING
  );
  PORT (
    clk, we : IN STD_LOGIC;
    adr : IN STD_LOGIC_VECTOR(ADDR - 1 DOWNTO 0);
    din : IN STD_LOGIC_VECTOR(DATA - 1 DOWNTO 0);
    dout : OUT STD_LOGIC_VECTOR(DATA - 1 DOWNTO 0)
  );
END;